`timescale 1ns / 1ps

module admin(
    
);


endmodule