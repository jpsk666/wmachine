`timescale 1ns / 1ps

module pre (
  input on,clk,rst,
  input p1,p2,p3,sign, //4个拨码开关，从右到左
  (* DONT_TOUCH = "1" *) 
  input r_pos,m_pos,u_pos,d_pos,//按键
  output reg isOn,  //按下按钮能否进入洗衣阶段
  output wire [7:0] led_r,  //数码管信号
  output [3:0] ena_r,  //数码管使能信号
  output wire [7:0] led_l,  //左数码管信号
  output [3:0] ena_l,  //左数码管使能信号
  output reg signed [11:0] bal,  //余额，最大999
  output reg [1:0] mode,  //模式 //有4个
  output reg [2:0] st_light  //接左边3小灯表示状态
);
reg [27:0] t;  //0.66秒计数
reg [3:0] n1, n2, n3, n0;  //1~3：个位至百位; 0:符号位
reg [3:0] n5, n6, n7, n8;  //1~3：个位至百位; 0:符号位
reg [29:0] alarm_t; //2.5s

parameter o = 1'b0;
parameter off = 4'hb;
parameter true = 1'b1;
wire next1;
assign next1 = ~(p1 | p2 | p3 | sign) & (n0 != 10);
//四个开关一个都不能上拨，且第一位不能是负数，才能下一阶段
reg [1:0] st = 1'b0;  //3种状态

wire m_pos,r_pos,u_pos,d_pos;
button bt(clk,bt,m_pos);
button bt_r(clk,bt_r,r_pos);
button bt_u(clk,bt_u,u_pos);
button bt_d(clk,bt_d,d_pos);

scan4 scanner (
    clk,
    n1,
    n2,
    n3,
    n0,
    ena_r,
    led_r
);
scan4 scanner2 (
    clk,
    n5,
    n6,
    n7,
    n8,
    ena_l,
    led_l
);

always @(*) begin  //小灯
  case (st)
    2'b00: begin //输入余额
      st_light <= 3'b001;
      isOn <= 0;
    end
    2'b01: begin //选择模式
      st_light <= 3'b010;
      isOn <= 0;
    end
    2'b10: begin //输入重量
      st_light <= 3'b100;
      case (mode)
        2'b01: begin
          if (n2 == 0 && d_pos) isOn <= 1;
          else isOn <= 0;
        end
        2'b10: begin
          if (n2 == 4'b000x && d_pos) isOn <= 1;
          else isOn <= 0;
        end
        default: begin
          if(d_pos) isOn <= 1;
        end
      endcase
    end
    default: begin
      st_light <= 3'b000;
      isOn <= 0;
    end
  endcase
end

always @(posedge clk, negedge rst) begin
  if (!rst) begin
    st <= 1'b0;
    {n1, n2, n3, n0} <= {o, o, o, o};
    {n5, n6, n7, n8} <= {off, off, off, off};
  end else begin
    if (on) begin
      case (st)  //状态判断
        2'b00: begin
          {n5, n6, n7, n8} <= {off, off, off, off};
          if (t >= 66000000) begin
            t <= 0;
            if (p1) begin  //拨上去时才加1,是否要写拨回去时的分支？
              if (n1 != 4'd9) n1 <= n1 + 1;
              else n1 <= 0;
            end else n1 <= n1;
            if (p2) begin
              if (n2 != 4'd9) n2 <= n2 + 1;
              else n2 <= 0;
            end else n2 <= n2;
            if (p3) begin
              if (n3 != 4'd9) n3 <= n3 + 1;
              else n3 <= 0;
            end else n3 <= n3;
            if (sign) begin
              if (n0 != 4'd10) n0 <= 4'd10;  //10代表负号
              else n0 <= 0;
            end else n0 <= n0;
          end else t <= t + 1;

          if (m_pos) begin  //如果按按钮就判断是否下一阶段
            if (next1) begin
              st <= 2'b01;
              n1 <= 0;  //可行，转化状态时直接赋值0
              {bal[4:1], bal[8:5], bal[12:9]} <= {n1, n2, n3};
              //可以这么做？
            end 
            else begin
              st <= 1'b0;
              {n0, n1, n2, n3} <= {o, o, o, o};
            end
          end else st <= 1'b0;
        end

        2'b01: begin
          {n5, n6, n7, n8} <= {off, off, off, off};
          {n2, n3, n0} <= {o, o, o};
          if (r_pos)
            if (n1 < 4'd3) n1 <= n1 + 1;
            else n1 <= 0;
          else n1 <= n1;

          if (u_pos) begin //开盖，进入下一状态
            st <= 2'b10;
            mode <= n1[1:0];//确定模式
            n8 <= n1;//放在最左侧显示
            {n0, n1, n2, n3} <= {o, o, o, o};
          end
        end
        2'b10: begin  //状态3
          //仍然是右按键增大
          if (r_pos) begin
            if (p1)//最右侧拨码开关上拨时表示十位数
              if (n2 > 4'd2)  //十位最多为20
                n2 <= 0;
              else n2 <= n2 + 1;
            else begin
              if (1 < 4'd9) n1 <= n1 + 1;
              else n1 <= 0;
            end
          end
          //确认输入
          if(m_pos)begin
            if(~isOn) begin
              case (mode)
              2'b00:begin //甩干
                if(n1 + n2*10<=) begin 
                  isOn<=1;
                end
              end
              2'b01:begin //小
                if(n1 + n2*10<=) begin 
                  isOn<=1;
                end
              end
              2'b10:begin //中
                if(n1 + n2*10<=) begin 
                  isOn<=1;
                end
              end
              2'b11:begin //大
                if(n1 + n2*10<=) begin 
                  isOn<=1;
                end
              end
              endcase
            end 
          end
        end
      endcase
    end
  end
end
endmodule

